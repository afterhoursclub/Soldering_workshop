.SUBCKT SN74HCS72 Data CLK CLR PRE Q Q_N VCC GND
XU6         11 PRE GND VCC GND BUFFER_0_0
XU5         12 CLR GND VCC GND BUFFER_0_0
XU10        Q_N 13 OE VCC GND BUFFER_0_0
XU9         Q 14 OE VCC GND BUFFER_0_0
XU8         16 15 CLK VCC GND BUFFER_0_0
XU1         17 Data CLKn VCC GND BUFFER_0_0
C2          13 GND 1P 
C1          18 GND 1P 
XU12        13 12 14 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU7         18 11 15 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU4         14 11 16 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
XU3         15 17 12 VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
R2          17 18 1K 
R1          16 13 1K 
XU2         CLKn VCC CLK VCC GND GATE_2INPUT_HC_2I_NAND_PP_ST_0
.ENDS


********************************************************************************
*                                 HCS_BUFFER
********************************************************************************

.SUBCKT BUFFER_0_0   Y A OEZ VCC AGND
XU1 Y A OEZ VCC AGND DRIVER_1INPUT_HC_1I_AND_TRISTATE_ST
.ENDS 

.SUBCKT DRIVER_1INPUT_HC_1I_AND_TRISTATE_ST Y A OEZ VCC AGND
XU1 Y A VCC OEZ VCC AGND LOGIC_GATE_2PIN_TRI_STATE_HC_1I_AND_TRISTATE_ST
.ENDS




*$
.SUBCKT LOGIC_GATE_2PIN_TRI_STATE_HC_1I_AND_TRISTATE_ST OUT A B OEZ VCC GND

.PARAM VCC_ABS_MAX = 7
.PARAM VCC_MAX = 6
.PARAM RA = 24000000000
.PARAM RB = 24000000000
.PARAM CA = 1E-08
.PARAM CB = 1E-08
.PARAM ROEZ = 5000
.PARAM COEZ = 3E-12
RA  A  GND {RA}
RB  B  GND {RB}
CA  A  GND {CA}
CB  B  GND {CB}
ROEZ OEZ GND {ROEZ}
COEZ OEZ GND {COEZ}
XUA NA A VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_ST
XUB NB B VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_ST
XUOEZ NOEZ OEZ VCC GND LOGIC_INPUT_HC_1I_AND_TRISTATE_ST
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_1I_AND_TRISTATE_ST
XOUTPD NOUTG NOUTTPD VCC GND TPD_HC_1I_AND_TRISTATE_ST
XUOUT NOUTTPD NOUT_INT NOEZ VCC GND LOGIC_TRI_STATE_OUTPUT_HC_1I_AND_TRISTATE_ST
XICC VCC GND NVIOUT LOGIC_ICC_HC_1I_AND_TRISTATE_ST
SICC VCC GND VCC GND SW1
* MONITOR OUTPUT CURRENT *
H1 NVIOUT GND VIOUT 1 
VIOUT NOUT_INT OUTSW 0 
SIOFF OUTSW OUT VCC GND SW2
DA2 GND A D1
DB2 GND B D1
DO2 GND OUT D1
DOE1 NOEZ VCC D1
DOE2 GND OEZ D1
RDA1 NA1 GND 100E6
SDA1 NA1 A VCC GND SW2
RDB1 NB1 GND 100E6
SDB1 NB1 B VCC GND SW2
SDO1 NO1 OUT VCC GND SW2
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60E6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10M ROFF = 100E6
.MODEL D1 D
.ENDS
*$
.SUBCKT LOGIC_INPUT_HC_1I_AND_TRISTATE_ST OUT IN VCC VEE
.PARAM STANDARD_INPUT_SELECT = 0

.PARAM SCHMITT_TRIGGER_INPUT_SELECT = 1
ESTD_THR VSTD_THR VEE TABLE {V(VCC,VEE)} =
+(1,0.5)
+(1.8,0.9)
+(2.5,1.25)
+(3.3,1.65)
+(5,2.5)
+(6,3)
ETRP_P VTRP_P VEE TABLE {V(VCC,VEE)} =
+(2,1.2)
+(4.5,2.5)
+(6,3.3)
ETRP_N VTRP_N VEE TABLE {V(VCC,VEE)} =
+(2,0.6)
+(4.5,1.6)
+(6,2)
EHYST VHYST VEE TABLE {V(VCC,VEE)} =
+(2,0.6)
+(4.5,0.9)
+(6,1.3)
ETRUE NTRUE VEE VALUE = {V(VCC,VEE)}
EFALSE NFALSE VEE VALUE = {0}
EBETA BETA VEE VALUE = {V(VHYST,VEE)/(V(NTRUE,VEE) - V(NFALSE,VEE) + V(VHYST,VEE))}
EFB NFB VEE VALUE = {(1 - V(BETA,VEE))*V(IN,VEE) + V(BETA,VEE)*V(CURR_OUT,VEE)}
*EFB NFB VEE VALUE = {(1 - V(BETA,VEE))*V(IN,VEE) + V(BETA,VEE)*V(OUT,VEE)}
EREF NREF VEE VALUE = {0.5*(1 - V(BETA,VEE))*(V(VTRP_P,VEE) + V(VTRP_N,VEE)) 
+ + 0.5*V(BETA,VEE)*(V(NTRUE,VEE) + V(NFALSE,VEE))}
EDIFF NDIFF VEE VALUE = {V(NFB,NREF)}
*ECOMP OUT VEE VALUE = {0.5*V(VCC,VEE)*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
ESWITCH VSWITCH VEE VALUE = {0.5*(-SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
ESWITCH1 VSWITCH1 VEE VALUE = {0.5*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
GCOMP VEE CURR_OUT VALUE = {SCHMITT_TRIGGER_INPUT_SELECT*0.5*V(VCC,VEE)*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
GSTD VEE CURR_OUT VALUE = {STANDARD_INPUT_SELECT*0.5*V(VCC,VEE)*(SGN(V(IN,VSTD_THR)) + ABS(SGN(V(IN,VSTD_THR))))}
ROUT CURR_OUT VEE 1
EMID MID VEE VALUE = {0.5*(V(VCC,VEE) + V(VEE))}
EARG NARG VEE VALUE = {V(CURR_OUT,VEE) - V(MID,VEE)}
EOUT OUT VEE VALUE = {0.5*(SGN(V(NARG,VEE)) + ABS(SGN(V(NARG,VEE) ) ) )}
*EOUT OUT VEE CURR_OUT VEE 1
.PARAM MAXICC = 0.0009
.PARAM VT = .7
.PARAM VCC_MIN = 2

EV_VT1 VTN VEE VALUE = { VT }
EV_VT2 VTP VEE VALUE = { V(VCC,VEE) - VT }

ETEST TEST VEE VALUE = {.9*V(VCC,VEE)}

EVTHDIFF VTH_DIFF VEE VALUE = {V(IN,VSTD_THR)}
EVTHPDIFF VTHP_DIFF VEE VALUE = {V(IN,VTRP_P)}
EVTHNDIFF VTHN_DIFF VEE VALUE = {V(IN,VTRP_N)}
EVTNDIFF VTN_DIFF VEE VALUE = { V(IN,VTN) }
EVTPDIFF VTP_DIFF VEE VALUE = { V(IN,VTP) }


GICCVA VCC VEE VALUE = { (-ABS(( (1+SGN(V(VTN_DIFF,VEE)) ) )/2 -1) * 2*MAXICC*((V(IN,VEE)-VT)/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH,VEE)}
GICCVB VCC VEE VALUE = { (ABS(( (1+SGN(V(VTHP_DIFF,VEE)) ) )/2 -1) * 2*MAXICC*((V(IN,VEE)-VT)/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH,VEE)}

GICCVC VCC VEE VALUE = { ( ABS(  (1+SGN(V(VTHN_DIFF,VEE)) ) )/2     * 2*MAXICC*((V(IN,VEE)-(V(VCC,VEE)-VT))/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH1,VEE)}
GICCVD VCC VEE VALUE = { (-ABS(  (1+SGN(V(VTP_DIFF,VEE)) ) )/2     * 2*MAXICC*((V(IN,VEE)-(V(VCC,VEE)-VT))/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH1,VEE)}

.ENDS
*$
.SUBCKT LOGIC_FUNCTION_2_HC_1I_AND_TRISTATE_ST A B OUT VCC VEE
GAND  VEE N1 VALUE = {V(A,VEE)*V(B,VEE)} 
RN1 N1 VEE 1 
EOUT OUT VEE N1 VEE 1 
.ENDS 
*$
.SUBCKT  TPD_HC_1I_AND_TRISTATE_ST IN OUT VCC VEE
.PARAM TPDELAY1 = 1N
.PARAM RS = 10K
.PARAM CS = {-TPDELAY1/(RS*LOG(0.5))}
*ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
+(2,5)
+(4.5,2)
+(6,1)
*R1 IN N1 {RS}
G1 IN N1 VALUE = {V(IN,N1)/(V(NTPDNORM,VEE)*RS)}
RZ IN N1 10G
C1 N1 VEE {CS}
E1 N2 VEE VALUE = {0.5*(1 + SGN(V(N1,VEE) - 0.5))}
EOUT OUT VEE N2 VEE 1
.ENDS
.SUBCKT LOGIC_TRI_STATE_OUTPUT_HC_1I_AND_TRISTATE_ST IN OUT OEZ VCC VEE
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(2,500)
+(4.5,50)
+(6,38.4)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(2,100)
+(4.5,42.5)
+(6,28.8)
EOEZ N2 VEE VALUE = {1-V(OEZ,VEE)}
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)*V(N2,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*V(N2,VEE)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS
*$
.SUBCKT LOGIC_ICC_HC_1I_AND_TRISTATE_ST VCC VEE VIOUT
.PARAM ICC = 2.5E-09
.PARAM VCC_MAX = 6
.PARAM VCC_MIN = 2
GICC VCC VEE VALUE = {ICC*0.5*(1 + SGN(V(VCC,VEE) - VCC_MIN))}
EGNDF GNDF 0 VALUE = {0.5*(V(VCC) + V(VEE))}
GOUTP VCC GNDF VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
GOUTN GNDF VEE VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
.ENDS
*$


********************************************************************************
*                                 NAND_FLIPFLOP
********************************************************************************

.SUBCKT GATE_2INPUT_HC_2I_NAND_PP_ST_0  Y A B VCC AGND
XU1 Y A B VCC AGND LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST
.ENDS


*$
.SUBCKT LOGIC_GATE_2PIN_OD_HC_2I_NAND_PP_ST OUT A B VCC GND
.PARAM VCC_ABS_MAX = 7
.PARAM VCC_MAX = 6
.PARAM RA = 240000000
.PARAM RB = 240000000
.PARAM CA = 5E-15
.PARAM CB = 5E-15
.PARAM ROEZ = 5000
.PARAM COEZ = 3E-12
RA  A  GND {RA}
RB  B  GND {RB}
CA  A  GND {CA}
CB  B  GND {CB}
XUA NA A VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUB NB B VCC GND LOGIC_INPUT_HC_2I_NAND_PP_ST
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_2I_NAND_PP_ST
XUOUT NOUTG NOUT_INT VCC GND LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST
XICC VCC GND NVIOUT LOGIC_ICC_HC_2I_NAND_PP_ST
SICC VCC GND VCC GND SW1
* MONITOR OUTPUT CURRENT *
H1 NVIOUT GND VIOUT 1 
VIOUT NOUT_INT OUTSW 0 
SIOFF OUTSW OUT VCC GND SW2
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60E6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10M ROFF = 100E6
.ENDS
*$

.SUBCKT LOGIC_INPUT_HC_2I_NAND_PP_ST OUT IN VCC VEE
ESTD_THR VSTD_THR VEE TABLE {V(VCC,VEE)} =
+(1,0.5)
+(6,3)
** OUTPUT VOLTAGES **
***********************************
**** STANDARD INPUT MODEL *********
*********************************** 
GSTD VEE CURR_OUT VALUE = {0.5*V(VCC,VEE)*(SGN(V(IN,VSTD_THR)) + ABS(SGN(V(IN,VSTD_THR))))}
ROUT CURR_OUT VEE 1
EMID MID VEE VALUE = {0.5*(V(VCC,VEE) + V(VEE))}
EARG NARG VEE VALUE = {V(CURR_OUT,VEE) - V(MID,VEE)}
EOUT OUT VEE VALUE = {0.5*(SGN(V(NARG,VEE)) + ABS(SGN(V(NARG,VEE) ) ) )}
*EOUT OUT VEE CURR_OUT VEE 1
.ENDS


*$
.SUBCKT LOGIC_FUNCTION_2_HC_2I_NAND_PP_ST A B OUT VCC VEE
GNAND VEE N1 VALUE = {(1 - V(A,VEE)*V(B,VEE))}
RN1 N1 VEE 1
EOUT OUT VEE N1 VEE 1
.ENDS


*$
.SUBCKT LOGIC_PP_OUTPUT_HC_2I_NAND_PP_ST IN OUT VCC VEE
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(2,1)
+(6,1)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(2,1)
+(6,1)
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS
*


.SUBCKT LOGIC_ICC_HC_2I_NAND_PP_ST VCC VEE VIOUT
.PARAM ICC = 2.5E-08
.PARAM VCC_MAX = 6
.PARAM VCC_MIN = 2
*GICC VCC VEE VALUE = {ICC*V(VCC,VEE)/VCC_MAX}
GICC VCC VEE VALUE = {ICC*0.5*(1 + SGN(V(VCC,VEE) - VCC_MIN))}
*
* FLOATING GROUND AT MID-RAIL
EGNDF GNDF 0 VALUE = {0.5*(V(VCC) + V(VEE))}
*
GOUTP VCC GNDF VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
GOUTN GNDF VEE VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
*
*GOUTP VCC GNDF VALUE = {IF(V(VIMON,GNDF) > 0, V(VIMON,GNDF),0)}
*GOUTN GNDF VEE VALUE = {IF(V(VIMON,GNDF) <= 0, V(VIMON,GNDF),0)}
.ENDS
*$
